module signExt #(
    parameters
) (
    port_list
);
    
endmodule